`timescale 1ns / 1ps
module CLA(
input [15:0] x,
input [15:0] y,
input cin,
output cout,
output [15:0] sum
    );

// P = x^y
// G = x&y
// Digital Design book expressions:
// Si = Pi ^^ Ci
// Ci+1 = Gi + PiCi 

// C1 = G0 + P0Cin
// C2 = G1 + P1(G0+P0Cin)
// C3 = G2 + P2(G1+(P1(G0+P0Cin)))
// C4 = G3 + P3(G2 + P2(G1+(P1(G0+P0Cin))))
wire [15:0] p,g,c;
assign p = x^y; 
assign g = x&y;
assign c[0] = cin;
assign c[1] = g[0] | (p[0]&cin);
assign c[2] = g[1] | (p[1]&(g[0] | (p[0]&cin)));
assign c[3] = g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))));
assign c[4] = g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))));
assign c[5] = g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))));
assign c[6] = g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))));
assign c[7] = g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))));
assign c[8] = g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))));
assign c[9] = g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))));
assign c[10] = g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))));
assign c[11] = g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))));
assign c[12] = g[11] | (p[11] & (g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))))));
assign c[13] = g[12] | (p[12] & (g[11] | (p[11] & (g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))))))));
assign c[14] = g[13] | (p[13] & (g[12] | (p[12] & (g[11] | (p[11] & (g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))))))))));
assign c[15] = g[14] | (p[14] &(g[13] | (p[13] & (g[12] | (p[12] & (g[11] | (p[11] & (g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))))))))))));
assign cout = g[15] | (p[15] & (g[14] | (p[14] &(g[13] | (p[13] & (g[12] | (p[12] & (g[11] | (p[11] & (g[10] | (p[10] & (g[9] | (p[9] & (g[8] | (p[8] & (g[7] | (p[7] & (g[6] | (p[6] & (g[5] | (p[5] & (g[4] | (p[4] & (g[3] | (p[3]& (g[2] | (p[2]&(g[1] | (p[1]&(g[0] | (p[0]&cin)))))))))))))))))))))))))))))));
 
assign sum = p^c;

endmodule
